`define CYCLE_TIME 50            

module TestBench;

reg                Clk;
reg                Start;
reg                Reset;
integer            i, outfile, counter;
integer            stall, flush;
parameter          num_cycles = 64;

always #(`CYCLE_TIME/2) Clk = ~Clk;    

CPU CPU(
    .clk_i  (Clk),
    .rst_i  (Reset)
);
  
initial begin
    $dumpfile("CPU.vcd");
    $dumpvars;
    counter = 0;
    stall = 0;
    flush = 0;
    
    // initialize instruction memory
    for(i=0; i<256; i=i+1) begin
        CPU.Instruction_Memory.memory[i] = 32'b0;
    end
    
    // initialize data memory
    for(i=0; i<32; i=i+1) begin
        CPU.Data_Memory.memory[i] = 32'b0;
    end    
        
    // Load instructions into instruction memory
    // Make sure you change back to "instruction.txt" before submission
    $readmemb("instruction.txt", CPU.Instruction_Memory.memory);
    
    // Open output file
    // Make sure you change back to "output.txt" before submission
    outfile = $fopen("output.txt") | 1;
    
    Clk = 0;
    Reset = 1;

    #(`CYCLE_TIME/8) 
    Reset = 0;

    #(`CYCLE_TIME/8) 
    Reset = 1;

    // [D-MemoryInitialization] DO NOT REMOVE THIS FLAG !!!
    CPU.Data_Memory.memory[0] = 5;
    CPU.Data_Memory.memory[1] = 6;
    CPU.Data_Memory.memory[2] = 10;
    CPU.Data_Memory.memory[3] = 18;
    CPU.Data_Memory.memory[4] = 29;

    CPU.Registers.register[24] = -24;
    CPU.Registers.register[25] = -25;
    CPU.Registers.register[26] = -26;
    CPU.Registers.register[27] = -27;
    CPU.Registers.register[28] = 56;
    CPU.Registers.register[29] = 58;
    CPU.Registers.register[30] = 60;
    CPU.Registers.register[31] = 62;

    // Pipeline Reg initialization
    CPU.ID_Pipeline_Reg.instr_out = 32'b0;
    CPU.ID_Pipeline_Reg.PC_out = 32'b0;

    CPU.EX_Pipeline_Reg.RegWrite_out = 1'b0;
    CPU.EX_Pipeline_Reg.MemtoReg_out = 1'b0;
    CPU.EX_Pipeline_Reg.MemRead_out = 1'b0;
    CPU.EX_Pipeline_Reg.MemWrite_out = 1'b0;
    CPU.EX_Pipeline_Reg.ALUOp_out = 2'b0;
    CPU.EX_Pipeline_Reg.ALUSrc_out = 1'b0;
    CPU.EX_Pipeline_Reg.data1_out = 32'b0;
    CPU.EX_Pipeline_Reg.data2_out = 32'b0;
    CPU.EX_Pipeline_Reg.immi_out = 32'b0;
    CPU.EX_Pipeline_Reg.funct_out = 10'b0;
    CPU.EX_Pipeline_Reg.Rs1_out = 5'b0;
    CPU.EX_Pipeline_Reg.Rs2_out = 5'b0;
    CPU.EX_Pipeline_Reg.Rd_out = 5'b0;

    CPU.MEM_Pipeline_Reg.RegWrite_out = 1'b0;
    CPU.MEM_Pipeline_Reg.MemtoReg_out = 1'b0;
    CPU.MEM_Pipeline_Reg.MemRead_out = 1'b0;
    CPU.MEM_Pipeline_Reg.MemWrite_out = 1'b0;
    CPU.MEM_Pipeline_Reg.ALU_result_out = 32'b0;
    CPU.MEM_Pipeline_Reg.data_2_out = 32'b0;
    CPU.MEM_Pipeline_Reg.Rd_out = 5'b0;

    CPU.WB_Pipeline_Reg.RegWrite_out = 1'b0;
    CPU.WB_Pipeline_Reg.MemtoReg_out = 1'b0;
    CPU.WB_Pipeline_Reg.data_ALU_out = 32'b0;
    CPU.WB_Pipeline_Reg.data_mem_out = 32'b0;
    CPU.WB_Pipeline_Reg.Rd_out = 5'b0;
    
    // Control Signal initialization
    CPU.Control.ALUOp = 2'b0;
    CPU.Control.ALUSrc = 1'b0;
    CPU.Control.RegWrite = 1'b0;
    CPU.Control.MemtoReg = 1'b0;
    CPU.Control.MemRead = 1'b0;
    CPU.Control.MemWrite = 1'b0;
    CPU.Control.Branch = 1'b0;

end
  
always@(posedge Clk) begin
    if(counter == num_cycles)    // stop after num_cycles cycles
        $finish;

    // put in your own signal to count stall and flush
    // if(CPU.Hazard_Detection.Stall_o == 1 && CPU.Control.Branch_o == 0)stall = stall + 1;
    // if(CPU.ID_FlushIF == 1)flush = flush + 1;
    if(CPU.Hazard_Detection_Unit.IF_ID_write == 0 && CPU.Control.Branch == 0)stall = stall + 1;
    if(CPU.ID_Pipeline_Reg.Flush == 1)flush = flush + 1;

    // print PC
    // DO NOT CHANGE THE OUTPUT FORMAT
    $fdisplay(outfile, "cycle = %d, Stall = %0d, Flush = %0d\nPC = %d", counter, stall, flush, CPU.PC.pc_o);
    
    // print Registers
    // DO NOT CHANGE THE OUTPUT FORMAT
    $fdisplay(outfile, "Registers");
    $fdisplay(outfile, "x0 = %d, x8  = %d, x16 = %d, x24 = %d", CPU.Registers.register[0], CPU.Registers.register[8] , CPU.Registers.register[16], CPU.Registers.register[24]);
    $fdisplay(outfile, "x1 = %d, x9  = %d, x17 = %d, x25 = %d", CPU.Registers.register[1], CPU.Registers.register[9] , CPU.Registers.register[17], CPU.Registers.register[25]);
    $fdisplay(outfile, "x2 = %d, x10 = %d, x18 = %d, x26 = %d", CPU.Registers.register[2], CPU.Registers.register[10], CPU.Registers.register[18], CPU.Registers.register[26]);
    $fdisplay(outfile, "x3 = %d, x11 = %d, x19 = %d, x27 = %d", CPU.Registers.register[3], CPU.Registers.register[11], CPU.Registers.register[19], CPU.Registers.register[27]);
    $fdisplay(outfile, "x4 = %d, x12 = %d, x20 = %d, x28 = %d", CPU.Registers.register[4], CPU.Registers.register[12], CPU.Registers.register[20], CPU.Registers.register[28]);
    $fdisplay(outfile, "x5 = %d, x13 = %d, x21 = %d, x29 = %d", CPU.Registers.register[5], CPU.Registers.register[13], CPU.Registers.register[21], CPU.Registers.register[29]);
    $fdisplay(outfile, "x6 = %d, x14 = %d, x22 = %d, x30 = %d", CPU.Registers.register[6], CPU.Registers.register[14], CPU.Registers.register[22], CPU.Registers.register[30]);
    $fdisplay(outfile, "x7 = %d, x15 = %d, x23 = %d, x31 = %d", CPU.Registers.register[7], CPU.Registers.register[15], CPU.Registers.register[23], CPU.Registers.register[31]);

    // print Data Memory
    // DO NOT CHANGE THE OUTPUT FORMAT
    $fdisplay(outfile, "Data Memory: 0x00 = %10d", CPU.Data_Memory.memory[0]);
    $fdisplay(outfile, "Data Memory: 0x04 = %10d", CPU.Data_Memory.memory[1]);
    $fdisplay(outfile, "Data Memory: 0x08 = %10d", CPU.Data_Memory.memory[2]);
    $fdisplay(outfile, "Data Memory: 0x0C = %10d", CPU.Data_Memory.memory[3]);
    $fdisplay(outfile, "Data Memory: 0x10 = %10d", CPU.Data_Memory.memory[4]);
    $fdisplay(outfile, "Data Memory: 0x14 = %10d", CPU.Data_Memory.memory[5]);
    $fdisplay(outfile, "Data Memory: 0x18 = %10d", CPU.Data_Memory.memory[6]);
    $fdisplay(outfile, "Data Memory: 0x1C = %10d", CPU.Data_Memory.memory[7]);

    $fdisplay(outfile, "\n");
    
    counter = counter + 1;
    
      
end

  
endmodule
